//-----------------------------------------------------------------------------
// Verilog 2001 (IEEE Std 1364-2001)
//-----------------------------------------------------------------------------
// Purpose  : ICG Cell
//------------------------------------------------------------------------------
// Process  : Intel
//------------------------------------------------------------------------------
//
// Author   : Kathleen Feng
// Date     : 18 October 2023
//------------------------------------------------------------------------------

module AhaClockGate (
    input   wire            TE,
    input   wire            E,
    input   wire            CP,
    output  wire            Q
);
    // Instantiate ICG cell here
    b15cilb01hn1n16x5 u_icg (
        .te                     (TE),
        .en                     (E),
        .clk                    (CP),
        .clkout                 (Q)
    );
endmodule
