module PCORNER
	(
	VSSPST, 
	VSS, 
	VDDPST, 
	VDD
	);
   inout VSSPST;
   inout VSS;
   inout VDDPST;
   inout VDD;
endmodule
