module Tbench;
  // ----------------------------------------------------------------------------
  // Debug and Trace
  // ----------------------------------------------------------------------------
  wire          nTRST;                     // Test reset
  wire          TMS;                       // Test Mode Select/SWDIN
  wire          TCK;                       // Test clock / SWCLK
  wire          TDI;                       // Test Data In
  wire          TDO;                       // Test Data Out

  // ----------------------------------------------------------------------------
  // UART
  // ----------------------------------------------------------------------------
  wire          uart0_txd;
  wire          uart0_rxd;
  wire          uart1_txd;
  wire          uart1_rxd;

  //-----------------------------------------
  // Clocks and reset
  //-----------------------------------------
  localparam MAIN_PERIOD    = 1.0;

  reg           master_clk;
  reg           po_reset_n;

  initial
  begin
    master_clk    = 1'b1;
  end

  always #(MAIN_PERIOD/2)  master_clk = ~master_clk;

  integer count;
  integer flag;
  integer start_time;
  integer start_time2;

  initial
  begin
    $set_toggle_region(Tbench);
    //$toggle_start();
    count = 0;
    flag = 0;
	start_time = 0;
    start_time2 = 0;
  end

  always@(posedge master_clk) begin
	
  if(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.stream_data_valid_g2f != 1'b0) begin
    if (count == 0) begin
      $toggle_start();
	  $display("count %d, start kernel", count);
	  start_time = $time;
    end
    if (count == 1) begin
  	  $toggle_stop();
      $toggle_report("run_1_kernel_plus_setup.saif", 1e-12,"Tbench");
	  $display("count %d, stop, time %d", count, $time - start_time);
  	  $toggle_reset();
    end
    count = count + 1;
  end
  

  if(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.pc_start_pulse != 1'b0) begin
    flag = 1;
    $toggle_start();
	$display("start reconfigure", count);
    start_time2 = $time;
  end

  if(flag && (Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.pcfg_g2f_interrupt_pulse != 1'b0)) begin
    flag = 0;
  	$toggle_stop();
    $toggle_report("reconfigure.saif", 1e-12,"Tbench");
	$display("stop, time %d", $time - start_time2);
  	$toggle_reset();
  end
  
  //if(Tbench.u_cmsdk_uart_capture_ard.reg_end_simulation == 1'b1) begin
  //	$toggle_stop();
  //    $toggle_report("conv3_3.saif", 1e-12,"Tbench");
  //end
  end

  initial  
  begin
    force Tbench.u_soc.pad_TLX_FWD_PAYLOAD_TDATA_HI = 24'b0;
    force Tbench.u_soc.pad_TLX_FWD_FLOW_TDATA = 2'b0;
    force Tbench.u_soc.pad_CGRA_JTAG_TDO = 1'b0;
    force Tbench.u_soc.pad_TPIU_TRACE_CLK = 1'b0;
    force Tbench.u_soc.pad_TPIU_TRACE_DATA = 1'b0;
    force Tbench.u_soc.pad_TPIU_TRACE_SWO = 1'b0;
    force Tbench.u_soc.pad_TLX_REV_PAYLOAD_TDATA_LO = 45'b0;
    force Tbench.u_soc.pad_TLX_REV_PAYLOAD_TDATA_HI = 35'b0;
    force Tbench.u_soc.pad_TLX_REV_FLOW_TDATA = 3'b0;
    force Tbench.u_soc.pad_TLX_FWD_PAYLOAD_TDATA_LO = 16'b0;
    force Tbench.u_soc.pad_TLX_FWD_CLK = 16'b0;
    force Tbench.u_soc.pad_LOOP_BACK = 16'b0;
    force Tbench.u_soc.IOPAD_left_LOOP_BACK_0.I = 16'b0;
    force Tbench.u_soc.IOPAD_left_TLX_FWD_CLK_0.I = 16'b0;
    force Tbench.u_soc.core.u_aha_platform_ctrl.CGRA_JTAG_RESETn = 1'b0;
    $deposit(Tbench.u_cmsdk_uart_capture_ard.reg_end_simulation, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.u_clk_selector_sys_clk.u_by1_clk_switch.clk_sel_reg.Q, 1'b0); 
    $deposit(Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.u_clk_selector_sys_clk.u_by1_clk_switch.clk_en_reg.Q, 1'b0); 
    $deposit(Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.u_clk_selector_sys_clk.u_by2_clk_switch.clk_sel_reg.Q, 1'b0); 
    $deposit(Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.u_clk_selector_sys_clk.u_by2_clk_switch.clk_en_reg.Q, 1'b0); 
    $deposit(Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.u_clk_selector_sys_clk.u_by4_clk_switch.clk_sel_reg.Q, 1'b0); 
    $deposit(Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.u_clk_selector_sys_clk.u_by4_clk_switch.clk_en_reg.Q, 1'b0); 
    $deposit(Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.u_clk_selector_sys_clk.u_by8_clk_switch.clk_sel_reg.Q, 1'b0); 
    $deposit(Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.u_clk_selector_sys_clk.u_by8_clk_switch.clk_en_reg.Q, 1'b0); 
    $deposit(Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.u_clk_selector_sys_clk.u_by16_clk_switch.clk_sel_reg.Q, 1'b0); 
    $deposit(Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.u_clk_selector_sys_clk.u_by16_clk_switch.clk_en_reg.Q, 1'b0); 
    $deposit(Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.u_clk_selector_sys_clk.u_by32_clk_switch.clk_sel_reg.Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.u_clk_selector_sys_clk.u_by32_clk_switch.clk_en_reg.Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0.axi_controller_axi_rvalid_reg.Q, 1'b0);

    // glb_tile[0] WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // glb_tile[0] CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // glb_tile[0] BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);


    // glb_tile[1]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);




    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);



    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);



    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);



    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);



    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);



    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);



    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);



    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);


    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);



    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);



    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);



    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);




    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);



    // glb_tile[0]
    // WEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_WEB_array_d1_reg_7 .Q, 1'b1);

    // CEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_CEB_array_d1_reg_7 .Q, 1'b1);

    // BWEB
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_0 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_1 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_2 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_3 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_4 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_5 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_6 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_7 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_8 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_9 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_10 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_11 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_12 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_13 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_14 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_15 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_16 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_17 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_18 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_19 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_20 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_21 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_22 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_23 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_24 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_25 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_26 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_27 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_28 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_29 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_30 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_31 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_32 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_33 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_34 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_35 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_36 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_37 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_38 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_39 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_40 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_41 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_42 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_43 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_44 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_45 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_46 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_47 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_48 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_49 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_50 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_51 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_52 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_53 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_54 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_55 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_56 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_57 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_58 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_59 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_60 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_61 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_62 .Q, 1'b1);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_BWEB_d1_reg_63 .Q, 1'b1);

    // A
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_A_to_mem_d1_reg_10 .Q, 1'b0);

    // D
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[0].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_0 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_1 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_2 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_3 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_4 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_5 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_6 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_7 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_8 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_9 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_10 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_11 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_12 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_13 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_14 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_15 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_16 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_17 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_18 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_19 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_20 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_21 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_22 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_23 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_24 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_25 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_26 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_27 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_28 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_29 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_30 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_31 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_32 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_33 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_34 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_35 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_36 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_37 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_38 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_39 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_40 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_41 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_42 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_43 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_44 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_45 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_46 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_47 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_48 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_49 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_50 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_51 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_52 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_53 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_54 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_55 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_56 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_57 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_58 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_59 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_60 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_61 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_62 .Q, 1'b0);
    $deposit(Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile .\glb_tile_int_glb_core_glb_bank_gen[1].bank_glb_bank_memory_glb_bank_sram_gen_D_d1_reg_63 .Q, 1'b0);



//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X00_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0A_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0C_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0D_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0E_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X01_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1A_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1C_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1D_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1E_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X02_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X04_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X05_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X06_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X08_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X09_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X10_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X11_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X12_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X14_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X15_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X16_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X18_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_PE.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X19_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0B_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X0F_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1B_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X1F_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X03_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X07_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X13_Y10,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y0A,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y0B,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y0C,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y0D,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y0E,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y0F,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y01,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y02,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y03,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y04,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y05,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y06,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y07,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y08,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y09,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/Tile_MemCore.sdf", Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0.Tile_X17_Y10,,,"MAXIMUM");
//
//$sdf_annotate("./inputs/gate_level/tile_array.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.Interconnect_inst0,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[0].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[1].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[2].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[3].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[4].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[5].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[6].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[7].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[8].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[9].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[10].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[11].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[12].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[13].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[14].glb_tile ,,,"MAXIMUM");
//$sdf_annotate("./inputs/gate_level/glb_tile.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0.\glb_tile_gen[15].glb_tile ,,,"MAXIMUM");
//
//$sdf_annotate("./inputs/gate_level/glb_top.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalBuffer_16_32_inst0$global_buffer_inst0,,,"MAXIMUM");
//
//$sdf_annotate("./inputs/gate_level/global_controller.sdf",Tbench.u_soc.core.u_aha_garnet.u_garnet.GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0);
//
//
//$sdf_annotate("inputs/gate_level/design.sdf",Tbench.u_soc,,"sdf_soc.log","MAXIMUM");
  end 






  initial
    begin
      po_reset_n   = 1'b0;
      #2000
      po_reset_n   = 1'b1;
    end

  //-----------------------------------------
  // AHASOC Integration
  //-----------------------------------------
  // TLX FWD Wires
  wire                                  tlx_fwd_clk;
  wire                                  tlx_fwd_payload_tvalid;
  wire                                  tlx_fwd_payload_tready;
  wire [(`TLX_FWD_DATA_LO_WIDTH-1):0]   tlx_fwd_payload_tdata_lo;
  wire [(39-`TLX_FWD_DATA_LO_WIDTH):0]  tlx_fwd_payload_tdata_hi;
  wire [39:0]                           tlx_fwd_payload_tdata;

  wire                                  tlx_fwd_flow_tvalid;
  wire                                  tlx_fwd_flow_tready;
  wire [1:0]                            tlx_fwd_flow_tdata;

  assign tlx_fwd_payload_tdata = {tlx_fwd_payload_tdata_hi, tlx_fwd_payload_tdata_lo};

  // TLX REV Wires
  wire                                  tlx_rev_payload_tvalid;
  wire                                  tlx_rev_payload_tready;
  wire [(`TLX_REV_DATA_LO_WIDTH-1):0]   tlx_rev_payload_tdata_lo;
  wire [(79-`TLX_REV_DATA_LO_WIDTH):0]  tlx_rev_payload_tdata_hi;
  wire [79:0]                           tlx_rev_payload_tdata;

  wire                                  tlx_rev_flow_tvalid;
  wire                                  tlx_rev_flow_tready;
  wire [2:0]                            tlx_rev_flow_tdata;

  wire tlx_rev_lane_0;
  wire [79:0] tlx_rev_payload_tdata_w;

  assign tlx_rev_payload_tdata_w  = {tlx_rev_payload_tdata[79:1], tlx_rev_lane_0};
  assign tlx_rev_payload_tdata_lo = tlx_rev_payload_tdata_w[(`TLX_REV_DATA_LO_WIDTH-1):0];
  assign tlx_rev_payload_tdata_hi = tlx_rev_payload_tdata_w[79:`TLX_REV_DATA_LO_WIDTH];

  GarnetSOC_pad_frame u_soc (
    .pad_jtag_intf_i_phy_tck        (1'b0),
    .pad_jtag_intf_i_phy_tdi        (1'b0),
    .pad_jtag_intf_i_phy_tdo        (),
    .pad_jtag_intf_i_phy_tms        (1'b0),
    .pad_jtag_intf_i_phy_trst_n     (1'b1),
    .pad_ext_rstb                   (1'b0),
    .pad_ext_dump_start             (1'b0),

    .pad_PORESETn                   (po_reset_n),
    .pad_DP_JTAG_TRSTn              (nTRST),
    .pad_CGRA_JTAG_TRSTn            (1'b1),

    .pad_MASTER_CLK                 (master_clk),
    .pad_DP_JTAG_TCK                (TCK),
    .pad_CGRA_JTAG_TCK              (1'b0),

    .pad_DP_JTAG_TDI                (TDI),
    .pad_DP_JTAG_TMS                (TMS),
    .pad_DP_JTAG_TDO                (TDO),

    .pad_CGRA_JTAG_TDI              (1'b0),
    .pad_CGRA_JTAG_TMS              (1'b0),
    .pad_CGRA_JTAG_TDO              (),

    .pad_TPIU_TRACE_DATA            (),
    .pad_TPIU_TRACE_SWO             (),
    .pad_TPIU_TRACE_CLK             (),

    .pad_UART0_RXD                  (uart0_rxd),
    .pad_UART0_TXD                  (uart0_txd),
    .pad_UART1_RXD                  (uart1_rxd),
    .pad_UART1_TXD                  (uart1_txd),

    // TLX FWD
    .pad_TLX_FWD_CLK                (tlx_fwd_clk),
    .pad_TLX_FWD_PAYLOAD_TVALID     (tlx_fwd_payload_tvalid),
    .pad_TLX_FWD_PAYLOAD_TREADY     (tlx_fwd_payload_tready),
    .pad_TLX_FWD_PAYLOAD_TDATA_LO   (tlx_fwd_payload_tdata_lo),
    .pad_TLX_FWD_PAYLOAD_TDATA_HI   (tlx_fwd_payload_tdata_hi),

    .pad_TLX_FWD_FLOW_TVALID        (tlx_fwd_flow_tvalid),
    .pad_TLX_FWD_FLOW_TREADY        (tlx_fwd_flow_tready),
    .pad_TLX_FWD_FLOW_TDATA         (tlx_fwd_flow_tdata),

    // TLX REV
    .pad_TLX_REV_CLK                (master_clk),

    .pad_TLX_REV_PAYLOAD_TVALID     (tlx_rev_payload_tvalid),
    .pad_TLX_REV_PAYLOAD_TREADY     (tlx_rev_payload_tready),
    .pad_TLX_REV_PAYLOAD_TDATA_LO   (tlx_rev_payload_tdata_lo),
    .pad_TLX_REV_PAYLOAD_TDATA_HI   (tlx_rev_payload_tdata_hi),

    .pad_TLX_REV_FLOW_TVALID        (tlx_rev_flow_tvalid),
    .pad_TLX_REV_FLOW_TREADY        (tlx_rev_flow_tready),
    .pad_TLX_REV_FLOW_TDATA         (tlx_rev_flow_tdata),

    // LoopBack
    .pad_LOOP_BACK_SELECT           (4'h0),
    .pad_LOOP_BACK                  ()
  );

  // TLX Master Domain
  tlx_mem u_tlx_m_dom (
    // FWD Link
    .tlx_fwd_clk                    (tlx_fwd_clk),
    .tlx_fwd_reset_n                (po_reset_n),

    .tlx_fwd_payload_tvalid         (tlx_fwd_payload_tvalid),
    .tlx_fwd_payload_tready         (tlx_fwd_payload_tready),
    .tlx_fwd_payload_tdata          (tlx_fwd_payload_tdata),

    .tlx_fwd_flow_tvalid            (tlx_fwd_flow_tvalid),
    .tlx_fwd_flow_tready            (tlx_fwd_flow_tready),
    .tlx_fwd_flow_tdata             (tlx_fwd_flow_tdata),

    // REV Link
    .tlx_rev_clk                    (master_clk),
    .tlx_rev_reset_n                (po_reset_n),

    .tlx_rev_payload_tvalid         (tlx_rev_payload_tvalid),
    .tlx_rev_payload_tready         (tlx_rev_payload_tready),
    .tlx_rev_payload_tdata          (tlx_rev_payload_tdata),

    .tlx_rev_flow_tvalid            (tlx_rev_flow_tvalid),
    .tlx_rev_flow_tready            (tlx_rev_flow_tready),
    .tlx_rev_flow_tdata             (tlx_rev_flow_tdata)
  );

  //-----------------------------------------
  // Pullup and pulldown
  //-----------------------------------------
  pullup(TDI);
  pullup(TMS);
  pullup(TCK);
  pullup(nTRST);
  pullup(TDO);

  pullup(uart0_rxd);
  pullup(uart1_rxd);

  //-----------------------------------------
  // max cycle set
  //-----------------------------------------
  int max_cycle;
  initial begin
    if ($value$plusargs("MAX_CYCLE=%0d", max_cycle)) begin
      repeat (max_cycle) @(posedge master_clk);
      $display("\n%0t\tERROR: The %0d cycles marker has passed!", $time, max_cycle);
      $finish(2);
    end
  end

  //-----------------------------------------
  // UART Loop Back
  //-----------------------------------------
  assign uart0_rxd  = uart0_txd;
  assign uart1_rxd  = uart1_txd;

  //-------------------------------------------
  // CXDT instantiation
  //-------------------------------------------
  CXDT #(.IMAGENAME ("./CXDT.bin"))
  u_cxdt(.CLK       (master_clk),
         .PORESETn  (po_reset_n),
         .TDO       (TDO),
         .TDI       (TDI),
         .nTRST     (nTRST),
         .SWCLKTCK  (TCK),
         .SWDIOTMS  (TMS)
  );

  //-----------------------------------------
  // UART0 Capture
  //-----------------------------------------
  cmsdk_uart_capture_ard u_cmsdk_uart_capture_ard (
    .RESETn              (po_reset_n),    // Power on reset
    .CLK                 (Tbench.u_soc.core.u_aha_platform_ctrl.u_clock_controller.UART0_CLK),      // Clock
    .RXD                 (uart0_txd),     // Received data
    .SIMULATIONEND       (),
    .DEBUG_TESTER_ENABLE (),
    .AUXCTRL             (),
    .SPI0                (),
    .SPI1                (),
    .I2C0                (),
    .I2C1                (),
    .UART0               (),
    .UART1               ()
  );

  assign uart0_rxd = uart0_txd;

  //-----------------------------------------
  // TLX Traning Capture
  //-----------------------------------------

  AhaTlxTrainingMonitor u_tlx_capture (
    .FWD_CLK            (tlx_fwd_clk),
    .FWD_RESETn         (po_reset_n),
    .REV_CLK            (master_clk),
    .REV_RESETn         (po_reset_n),
    .OE                 (Tbench.u_soc.core.u_aha_tlx.u_aha_tlx_ctrl.l2h_LANE_ENABLE_REG_LANE0_r),
    .FWD_DATA_IN        (tlx_fwd_payload_tdata[0]),
    .REV_DATA_IN        (tlx_rev_payload_tdata[0]),
    .REV_DATA_OUT       (tlx_rev_lane_0)
  );

  //-----------------------------------------
  // VCD Dump
  //-----------------------------------------
  // dumping trn file can speed up
  initial begin
    if ($test$plusargs("VCD_ON")) begin
      //$recordfile("dump.trn");
      //$recordvars(Tbench);
      $vcdplusfile("dump.vpd");
      $vcdpluson;
    end
  end

endmodule
