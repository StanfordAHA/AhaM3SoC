module PCORNER (
    input wire RTE
);
    wire unused = RTE;
endmodule
